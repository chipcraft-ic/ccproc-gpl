// +FHDR------------------------------------------------------------------------
//
// Copyright (c) 2017 ChipCraft Sp. z o.o. All rights reserved
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, version 2.
//
// This program is distributed in the hope that it will be useful, but
// WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program. If not, see <http://www.gnu.org/licenses/>
//
// -----------------------------------------------------------------------------
// Author    : Krzysztof Marcinek
// -----------------------------------------------------------------------------
// $Date: 2017-03-30 21:39:22 +0200 (Thu, 30 Mar 2017) $
// $Revision: 21 $
// -FHDR------------------------------------------------------------------------

`ifndef __DEBUG_DEFINE__
`define __DEBUG_DEFINE__

`define DUMP_BLOCK_DEF 32'd26

`endif // __DEBUG_DEFINE__


// +FHDR------------------------------------------------------------------------
//
// Copyright (c) 2017 ChipCraft Sp. z o.o. All rights reserved
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, version 2.
//
// This program is distributed in the hope that it will be useful, but
// WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program. If not, see <http://www.gnu.org/licenses/>
//
// -----------------------------------------------------------------------------
// File Name : add.v
// Author    : Krzysztof Marcinek
// -----------------------------------------------------------------------------
// $Date: 2019-03-15 10:27:52 +0100 (Fri, 15 Mar 2019) $
// $Revision: 431 $
// -FHDR------------------------------------------------------------------------

`include "timescale.inc"
`include "define.vh"



// -----------------------------------------------------------------------------
// adder module with carry input
// -----------------------------------------------------------------------------

module addcin_module(a, b, cin, q);

// -----------------------------------------------------------------------------
// parameters
// -----------------------------------------------------------------------------

parameter [31:0] WIDTH = 32'd32;

// -----------------------------------------------------------------------------
// ports
// -----------------------------------------------------------------------------

input wire      [WIDTH-1:0]     a;
input wire      [WIDTH-1:0]     b;
input wire                      cin;
output wire     [WIDTH-1:0]     q;

// -----------------------------------------------------------------------------
// assign output
// -----------------------------------------------------------------------------

assign q = a + b + cin;

endmodule



// -----------------------------------------------------------------------------
// adder module with carry input and enable
// -----------------------------------------------------------------------------

module addcinen_module(a, b, cin, q, en);

// -----------------------------------------------------------------------------
// parameters
// -----------------------------------------------------------------------------

parameter [31:0] WIDTH = 32'd32;
parameter [31:0] OPIS  = 32'd32;

// -----------------------------------------------------------------------------
// ports
// -----------------------------------------------------------------------------

input wire      [WIDTH-1:0]     a;
input wire      [WIDTH-1:0]     b;
input wire                      cin;
input wire                      en;
output reg      [WIDTH-1:0]     q;

generate

// -----------------------------------------------------------------------------
// operand isolation
// -----------------------------------------------------------------------------

if (OPIS == 1) begin
    wire    [WIDTH-1:0]     isol_a;
    wire    [WIDTH-1:0]     isol_b;
    wire                    isol_cin;
    assign  isol_a     = a & {WIDTH{en}};
    assign  isol_b     = b & {WIDTH{en}};
    assign  isol_cin   = cin & en;
    always @(*)
    begin
        q = isol_a + isol_b + {{WIDTH-1{1'b0}},isol_cin};
    end
end

// -----------------------------------------------------------------------------
// without operand isolation
// -----------------------------------------------------------------------------

else begin
    always @(*)
    begin
        q = a + b + {{WIDTH-1{1'b0}},cin};
    end
end
endgenerate

endmodule



// -----------------------------------------------------------------------------
// adder module with carry out
// -----------------------------------------------------------------------------

module addcout_module(a, b, cout, q);

// -----------------------------------------------------------------------------
// parameters
// -----------------------------------------------------------------------------

parameter [31:0] WIDTH = 32'd32;

// -----------------------------------------------------------------------------
// ports
// -----------------------------------------------------------------------------

input wire      [WIDTH-1:0]     a;
input wire      [WIDTH-1:0]     b;
output wire                     cout;
output wire     [WIDTH-1:0]     q;

// -----------------------------------------------------------------------------
// assign output
// -----------------------------------------------------------------------------

assign {cout,q} = a + b;

endmodule



// -----------------------------------------------------------------------------
// adder module
// -----------------------------------------------------------------------------

module add_module(a, b, q);

// -----------------------------------------------------------------------------
// parameters
// -----------------------------------------------------------------------------

parameter [31:0] WIDTH = 32'd32;

// -----------------------------------------------------------------------------
// ports
// -----------------------------------------------------------------------------

input wire      [WIDTH-1:0]     a;
input wire      [WIDTH-1:0]     b;
output wire     [WIDTH-1:0]     q;

// -----------------------------------------------------------------------------
// assign output
// -----------------------------------------------------------------------------

assign q = a + b;

endmodule



// -----------------------------------------------------------------------------
// adder module with enable
// -----------------------------------------------------------------------------

module adden_module(a, b, en, q);

// -----------------------------------------------------------------------------
// parameters
// -----------------------------------------------------------------------------

parameter [31:0] WIDTH = 32'd32;
parameter [31:0] OPIS  = 32'd32;

// -----------------------------------------------------------------------------
// ports
// -----------------------------------------------------------------------------

input wire      [WIDTH-1:0]     a;
input wire      [WIDTH-1:0]     b;
input wire                      en;
output reg      [WIDTH-1:0]     q;

generate

// -----------------------------------------------------------------------------
// operand isolation
// -----------------------------------------------------------------------------

if (OPIS == 1) begin
    wire    [WIDTH-1:0]    isol_a;
    wire    [WIDTH-1:0]    isol_b;
    assign  isol_a = a & {WIDTH{en}};
    assign  isol_b = b & {WIDTH{en}};
    always @(*)
    begin
        q = isol_a + isol_b;
    end
end

// -----------------------------------------------------------------------------
// without operand isolation
// -----------------------------------------------------------------------------

else begin
    always @(*)
    begin
        q = a + b;
    end
end
endgenerate

endmodule



// -----------------------------------------------------------------------------
// adder module with carry out and enable
// -----------------------------------------------------------------------------

module addencout_module(a, b, en, q, cout);

// -----------------------------------------------------------------------------
// parameters
// -----------------------------------------------------------------------------

parameter [31:0] WIDTH = 32'd32;
parameter [31:0] OPIS  = 32'd32;

// -----------------------------------------------------------------------------
// ports
// -----------------------------------------------------------------------------

input wire  [WIDTH-1:0] a;
input wire  [WIDTH-1:0] b;
input wire              en;
output reg              cout;
output reg  [WIDTH-1:0] q;

generate

// -----------------------------------------------------------------------------
// opernad isolation
// -----------------------------------------------------------------------------

if (OPIS == 1) begin
    wire    [WIDTH-1:0] isol_a;
    wire    [WIDTH-1:0] isol_b;
    assign  isol_a = a & {WIDTH{en}};
    assign  isol_b = b & {WIDTH{en}};
    always @(*)
    begin
        {cout,q} = isol_a + isol_b;
    end
end

// -----------------------------------------------------------------------------
// without opernad isolation
// -----------------------------------------------------------------------------

else begin
    always @(*)
    begin
        {cout,q} = a + b;
    end
end
endgenerate

endmodule
